module constants

pub enum Response {
    argon2_ok = 0
argon_2_output_ptr_null_1 = -1

argon_2_output_too_short_2 = -2
argon_2_output_too_long_3 = -3

argon_2_pwd_too_short_4 = -4
argon_2_pwd_too_long_5 = -5

argon_2_salt_too_short_6 = -6
argon_2_salt_too_long_7 = -7

argon_2_ad_too_short_8 = -8
argon_2_ad_too_long_9 = -9

argon_2_secret_too_short_10 = -10
argon_2_secret_too_long_11 = -11

argon_2_time_too_small_12 = -12
argon_2_time_too_large_13 = -13

argon_2_memory_too_little_14 = -14
argon_2_memory_too_much_15 = -15

argon_2_lanes_too_few_16 = -16
argon_2_lanes_too_many_17 = -17

argon_2_pwd_ptr_mismatch_18 = -18
argon_2_salt_ptr_mismatch_19 = -19
argon_2_secret_ptr_mismatch_20 = -20
argon_2_ad_ptr_mismatch_21 = -21

argon_2_memory_allocation_error_22 = -22

argon_2_free_memory_cbk_null_23 = -23
argon_2_allocate_memory_cbk_null_24 = -24

argon_2_incorrect_parameter_25 = -25
argon_2_incorrect_type_26 = -26

argon_2_out_ptr_mismatch_27 = -27

argon_2_threads_too_few_28 = -28
argon_2_threads_too_many_29 = -29

argon_2_missing_args_30 = -30

argon_2_encoding_fail_31 = -31

argon_2_decoding_fail_32 = -32

argon_2_thread_fail_33 = -33

argon_2_decoding_length_fail_34 = -34

argon_2_verify_mismatch_35 = -35

    
	}