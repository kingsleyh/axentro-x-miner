module argon2

#flag -I @VROOT/c
#flag @VROOT/c/

#include "include/argon2.h"

